magic
tech sky130A
magscale 1 2
timestamp 1679269954
<< error_p >>
rect -29 522 29 528
rect -29 488 -17 522
rect -29 482 29 488
rect -29 -488 29 -482
rect -29 -522 -17 -488
rect -29 -528 29 -522
<< nmos >>
rect -15 -450 15 450
<< ndiff >>
rect -73 438 -15 450
rect -73 -438 -61 438
rect -27 -438 -15 438
rect -73 -450 -15 -438
rect 15 438 73 450
rect 15 -438 27 438
rect 61 -438 73 438
rect 15 -450 73 -438
<< ndiffc >>
rect -61 -438 -27 438
rect 27 -438 61 438
<< poly >>
rect -33 522 33 538
rect -33 488 -17 522
rect 17 488 33 522
rect -33 472 33 488
rect -15 450 15 472
rect -15 -472 15 -450
rect -33 -488 33 -472
rect -33 -522 -17 -488
rect 17 -522 33 -488
rect -33 -538 33 -522
<< polycont >>
rect -17 488 17 522
rect -17 -522 17 -488
<< locali >>
rect -33 488 -17 522
rect 17 488 33 522
rect -61 438 -27 454
rect -61 -454 -27 -438
rect 27 438 61 454
rect 27 -454 61 -438
rect -33 -522 -17 -488
rect 17 -522 33 -488
<< viali >>
rect -17 488 17 522
rect -61 -438 -27 438
rect 27 -438 61 438
rect -17 -522 17 -488
<< metal1 >>
rect -29 522 29 528
rect -29 488 -17 522
rect 17 488 29 522
rect -29 482 29 488
rect -67 438 -21 450
rect -67 -438 -61 438
rect -27 -438 -21 438
rect -67 -450 -21 -438
rect 21 438 67 450
rect 21 -438 27 438
rect 61 -438 67 438
rect 21 -450 67 -438
rect -29 -488 29 -482
rect -29 -522 -17 -488
rect 17 -522 29 -488
rect -29 -528 29 -522
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
