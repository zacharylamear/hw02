magic
tech sky130A
magscale 1 2
timestamp 1679269954
<< error_p >>
rect -29 2631 29 2637
rect -29 2597 -17 2631
rect -29 2591 29 2597
rect -29 -2597 29 -2591
rect -29 -2631 -17 -2597
rect -29 -2637 29 -2631
<< nwell >>
rect -109 -2650 109 2650
<< pmos >>
rect -15 -2550 15 2550
<< pdiff >>
rect -73 2538 -15 2550
rect -73 -2538 -61 2538
rect -27 -2538 -15 2538
rect -73 -2550 -15 -2538
rect 15 2538 73 2550
rect 15 -2538 27 2538
rect 61 -2538 73 2538
rect 15 -2550 73 -2538
<< pdiffc >>
rect -61 -2538 -27 2538
rect 27 -2538 61 2538
<< poly >>
rect -33 2631 33 2647
rect -33 2597 -17 2631
rect 17 2597 33 2631
rect -33 2581 33 2597
rect -15 2550 15 2581
rect -15 -2581 15 -2550
rect -33 -2597 33 -2581
rect -33 -2631 -17 -2597
rect 17 -2631 33 -2597
rect -33 -2647 33 -2631
<< polycont >>
rect -17 2597 17 2631
rect -17 -2631 17 -2597
<< locali >>
rect -33 2597 -17 2631
rect 17 2597 33 2631
rect -61 2538 -27 2554
rect -61 -2554 -27 -2538
rect 27 2538 61 2554
rect 27 -2554 61 -2538
rect -33 -2631 -17 -2597
rect 17 -2631 33 -2597
<< viali >>
rect -17 2597 17 2631
rect -61 -2538 -27 2538
rect 27 -2538 61 2538
rect -17 -2631 17 -2597
<< metal1 >>
rect -29 2631 29 2637
rect -29 2597 -17 2631
rect 17 2597 29 2631
rect -29 2591 29 2597
rect -67 2538 -21 2550
rect -67 -2538 -61 2538
rect -27 -2538 -21 2538
rect -67 -2550 -21 -2538
rect 21 2538 67 2550
rect 21 -2538 27 2538
rect 61 -2538 67 2538
rect 21 -2550 67 -2538
rect -29 -2597 29 -2591
rect -29 -2631 -17 -2597
rect 17 -2631 29 -2597
rect -29 -2637 29 -2631
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 25.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
