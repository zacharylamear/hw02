magic
tech sky130A
magscale 1 2
timestamp 1679318755
<< nwell >>
rect 630 2404 1152 2450
rect 630 2402 1156 2404
rect 796 2328 1156 2402
rect 794 2294 1156 2328
rect 790 2280 1156 2294
rect 790 2218 1134 2280
rect 1320 2274 1772 2446
<< pwell >>
rect 260 642 1332 1340
rect 260 168 1786 642
rect 256 -40 1786 168
rect 256 -64 656 -40
rect 694 -156 1786 -40
rect 694 -548 1288 -156
<< psubdiff >>
rect 786 -322 1186 -292
rect 786 -484 828 -322
rect 1140 -484 1186 -322
rect 786 -512 1186 -484
<< nsubdiff >>
rect 838 2378 1068 2404
rect 838 2294 862 2378
rect 1040 2294 1068 2378
rect 838 2268 1068 2294
<< psubdiffcont >>
rect 828 -484 1140 -322
<< nsubdiffcont >>
rect 862 2294 1040 2378
<< locali >>
rect 850 2402 886 2404
rect 850 2392 1064 2402
rect 850 2382 1068 2392
rect 850 2292 862 2382
rect 1044 2292 1068 2382
rect 850 2284 1068 2292
rect 850 2278 1064 2284
rect 850 2274 886 2278
rect 792 -320 1182 -296
rect 792 -482 818 -320
rect 1148 -482 1182 -320
rect 792 -484 828 -482
rect 1140 -484 1182 -482
rect 792 -510 1182 -484
<< viali >>
rect 862 2378 1044 2382
rect 862 2294 1040 2378
rect 1040 2294 1044 2378
rect 862 2292 1044 2294
rect 818 -322 1148 -320
rect 818 -482 828 -322
rect 828 -482 1140 -322
rect 1140 -482 1148 -322
<< metal1 >>
rect 1142 2596 1844 2598
rect 308 2452 772 2522
rect 1098 2456 1844 2596
rect 312 850 412 2452
rect 722 2390 768 2452
rect 1042 2402 1070 2404
rect 850 2390 1070 2402
rect 714 2382 1070 2390
rect 714 2292 862 2382
rect 1044 2380 1070 2382
rect 1098 2396 1202 2456
rect 1098 2380 1218 2396
rect 1044 2292 1218 2380
rect 714 2278 1218 2292
rect 714 2250 876 2278
rect 1034 2242 1218 2278
rect 538 1424 660 1668
rect 1260 1584 1584 1730
rect 910 1424 1278 1448
rect 490 1354 1278 1424
rect 490 1336 700 1354
rect 490 934 646 1336
rect 1432 932 1572 1584
rect 1886 936 2186 1212
rect 312 816 422 850
rect 314 630 422 816
rect 1234 746 1572 932
rect 1234 640 2016 746
rect 1234 630 1572 640
rect 314 540 490 630
rect 1234 618 1470 630
rect 382 320 490 540
rect 2088 538 2186 936
rect 1034 530 1176 532
rect 908 524 1176 530
rect 698 408 1176 524
rect 698 406 1070 408
rect 698 390 928 406
rect 156 206 322 306
rect 400 284 524 320
rect 380 224 524 284
rect 632 282 712 346
rect 854 278 928 390
rect 1694 386 2186 538
rect 1168 312 1242 380
rect 974 282 1140 286
rect 1274 282 1640 286
rect 126 164 252 206
rect 296 194 322 206
rect 126 -8 250 164
rect 400 158 524 224
rect 974 274 1640 282
rect 974 202 1338 274
rect 1520 202 1640 274
rect 974 186 1640 202
rect 312 146 858 158
rect 1110 146 1342 150
rect 312 78 1342 146
rect 958 74 1342 78
rect 126 -36 478 -8
rect 126 -172 160 -36
rect 128 -218 160 -172
rect 452 -120 478 -36
rect 1110 -42 1342 74
rect 1108 -50 1568 -42
rect 452 -218 890 -120
rect 1108 -144 1738 -50
rect 128 -256 890 -218
rect 364 -292 890 -256
rect 364 -320 1190 -292
rect 364 -432 818 -320
rect 790 -482 818 -432
rect 1148 -482 1190 -320
rect 790 -524 1190 -482
<< via1 >>
rect 1338 202 1520 274
rect 160 -218 452 -36
<< metal2 >>
rect 1302 274 1540 294
rect 1302 220 1338 274
rect 1216 202 1338 220
rect 1520 202 1540 274
rect 1216 180 1540 202
rect 130 -12 278 -10
rect 1216 -12 1396 180
rect 130 -36 1396 -12
rect 130 -218 160 -36
rect 452 -218 1396 -36
rect 130 -254 1396 -218
rect 1216 -256 1396 -254
use sky130_fd_pr__nfet_01v8_4WPVHQ  XM1
timestamp 1679278092
transform 1 0 953 0 1 243
box -73 -157 73 157
use sky130_fd_pr__pfet_01v8_LJPZDL  XM2
timestamp 1679278092
transform 1 0 1239 0 1 1898
box -109 -514 109 548
use sky130_fd_pr__nfet_01v8_FN4ZCM  XM4
timestamp 1679278092
transform 1 0 1203 0 1 829
box -73 -507 73 507
use sky130_fd_pr__pfet_01v8_27MD4L  XM7
timestamp 1679278092
transform 1 0 1863 0 1 3290
box -109 -2614 109 2648
use sky130_fd_pr__nfet_01v8_AT4ZK9  XM8
timestamp 1679278092
transform 1 0 1665 0 1 249
box -73 -357 73 357
use sky130_fd_pr__nfet_01v8_4WPVHQ  sky130_fd_pr__nfet_01v8_4WPVHQ_0
timestamp 1679278092
transform 1 0 353 0 1 255
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_FN4ZCM  sky130_fd_pr__nfet_01v8_FN4ZCM_0
timestamp 1679278092
transform 1 0 671 0 1 797
box -73 -507 73 507
use sky130_fd_pr__pfet_01v8_LJPZDL  sky130_fd_pr__pfet_01v8_LJPZDL_0
timestamp 1679278092
transform 1 0 687 0 1 1876
box -109 -514 109 548
<< labels >>
rlabel pwell 630 284 710 306 1 in_p
port 1 n
rlabel metal1 632 284 712 306 1 in_p
port 1 n
rlabel metal1 1052 2268 1118 2366 1 VDD
port 2 n
rlabel metal1 2054 990 2144 1110 1 diff_out
port 3 n
rlabel metal1 1172 314 1240 336 1 in_n
port 4 n
rlabel metal1 588 -400 772 -240 1 VSS
port 5 n
<< end >>
