magic
tech sky130A
magscale 1 2
timestamp 1679278092
<< error_p >>
rect -29 -461 29 -455
rect -29 -495 -17 -461
rect -29 -501 29 -495
<< nwell >>
rect -109 -514 109 548
<< pmos >>
rect -15 -414 15 486
<< pdiff >>
rect -73 474 -15 486
rect -73 -402 -61 474
rect -27 -402 -15 474
rect -73 -414 -15 -402
rect 15 474 73 486
rect 15 -402 27 474
rect 61 -402 73 474
rect 15 -414 73 -402
<< pdiffc >>
rect -61 -402 -27 474
rect 27 -402 61 474
<< poly >>
rect -15 486 15 512
rect -15 -445 15 -414
rect -33 -461 33 -445
rect -33 -495 -17 -461
rect 17 -495 33 -461
rect -33 -511 33 -495
<< polycont >>
rect -17 -495 17 -461
<< locali >>
rect -61 474 -27 490
rect -61 -418 -27 -402
rect 27 474 61 490
rect 27 -418 61 -402
rect -33 -495 -17 -461
rect 17 -495 33 -461
<< viali >>
rect -61 -402 -27 474
rect 27 -402 61 474
rect -17 -495 17 -461
<< metal1 >>
rect -67 474 -21 486
rect -67 -402 -61 474
rect -27 -402 -21 474
rect -67 -414 -21 -402
rect 21 474 67 486
rect 21 -402 27 474
rect 61 -402 67 474
rect 21 -414 67 -402
rect -29 -461 29 -455
rect -29 -495 -17 -461
rect 17 -495 29 -461
rect -29 -501 29 -495
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
