magic
tech sky130A
magscale 1 2
timestamp 1679278092
<< error_p >>
rect -29 -457 29 -451
rect -29 -491 -17 -457
rect -29 -497 29 -491
<< nmos >>
rect -15 -419 15 481
<< ndiff >>
rect -73 469 -15 481
rect -73 -407 -61 469
rect -27 -407 -15 469
rect -73 -419 -15 -407
rect 15 469 73 481
rect 15 -407 27 469
rect 61 -407 73 469
rect 15 -419 73 -407
<< ndiffc >>
rect -61 -407 -27 469
rect 27 -407 61 469
<< poly >>
rect -15 481 15 507
rect -15 -441 15 -419
rect -33 -457 33 -441
rect -33 -491 -17 -457
rect 17 -491 33 -457
rect -33 -507 33 -491
<< polycont >>
rect -17 -491 17 -457
<< locali >>
rect -61 469 -27 485
rect -61 -423 -27 -407
rect 27 469 61 485
rect 27 -423 61 -407
rect -33 -491 -17 -457
rect 17 -491 33 -457
<< viali >>
rect -61 -407 -27 469
rect 27 -407 61 469
rect -17 -491 17 -457
<< metal1 >>
rect -67 469 -21 481
rect -67 -407 -61 469
rect -27 -407 -21 469
rect -67 -419 -21 -407
rect 21 469 67 481
rect 21 -407 27 469
rect 61 -407 67 469
rect 21 -419 67 -407
rect -29 -457 29 -451
rect -29 -491 -17 -457
rect 17 -491 29 -457
rect -29 -497 29 -491
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
